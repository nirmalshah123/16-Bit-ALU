entity ALU_16_bit is

port (s0,s1 : in bit);		--S0,S1 are the control pins

end ALU_16_bit;

architecture M of ALU_16_bit is
begin
end M;
