entity ALU_16_bit is
port (A : in bit);
end ALU_16_bit;

architecture ALU of ALU_16_bit is
begin
end ALU;